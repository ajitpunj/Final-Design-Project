// mysystem.v

// Generated using ACDS version 13.1 162 at 2015.05.20.15:11:48

`timescale 1 ps / 1 ps
module mysystem (
		output wire [12:0] memory_mem_a,              //              memory.mem_a
		output wire [2:0]  memory_mem_ba,             //                    .mem_ba
		output wire        memory_mem_ck,             //                    .mem_ck
		output wire        memory_mem_ck_n,           //                    .mem_ck_n
		output wire        memory_mem_cke,            //                    .mem_cke
		output wire        memory_mem_cs_n,           //                    .mem_cs_n
		output wire        memory_mem_ras_n,          //                    .mem_ras_n
		output wire        memory_mem_cas_n,          //                    .mem_cas_n
		output wire        memory_mem_we_n,           //                    .mem_we_n
		output wire        memory_mem_reset_n,        //                    .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,             //                    .mem_dq
		inout  wire        memory_mem_dqs,            //                    .mem_dqs
		inout  wire        memory_mem_dqs_n,          //                    .mem_dqs_n
		output wire        memory_mem_odt,            //                    .mem_odt
		output wire        memory_mem_dm,             //                    .mem_dm
		input  wire        memory_oct_rzqin,          //                    .oct_rzqin
		output wire        hps_read_export,           //            hps_read.export
		output wire        vga_clk_clk,               //             vga_clk.clk
		output wire        d5m_clk_clk,               //             d5m_clk.clk
		output wire        dram_clk_clk,              //            dram_clk.clk
		output wire        sdram_clk_clk,             //           sdram_clk.clk
		input  wire        system_pll_0_reset_reset,  //  system_pll_0_reset.reset
		input  wire        system_pll_0_refclk_clk,   // system_pll_0_refclk.clk
		input  wire        sdram_clk_ref_clk_clk,     //   sdram_clk_ref_clk.clk
		input  wire        sdram_clk_ref_reset_reset, // sdram_clk_ref_reset.reset
		output wire        capture_start_export,      //       capture_start.export
		input  wire [15:0] sdram_hps_data1_export,    //     sdram_hps_data1.export
		input  wire [15:0] sdram_hps_data2_export,    //     sdram_hps_data2.export
		output wire [15:0] hps_vga_data1_export,      //       hps_vga_data1.export
		output wire [15:0] hps_vga_data2_export,      //       hps_vga_data2.export
		output wire        sdramclock_export,         //          sdramclock.export
		output wire        sdram_start_export,        //         sdram_start.export
		output wire        fifowe_export,             //              fifowe.export
		input  wire [9:0]  binary_export,             //              binary.export
		output wire [7:0]  greyparameter_export,      //       greyparameter.export
		input  wire        vgaclock_export,           //            vgaclock.export
		output wire        vgabinary_export,          //           vgabinary.export
		input  wire        vgaread_export,            //             vgaread.export
		input  wire [9:0]  topedge_export,            //             topedge.export
		output wire        hwreset_export,            //             hwreset.export
		input  wire        lval_export                //                lval.export
	);

	wire          sdram_clk_sdram_clk_clk;                                   // sdram_clk:sdram_clk_clk -> [FIFOWe:clk, Lval:clk, Onchip_SRAM:clk, Sdram_start:clk, arm_a9_hps:f2h_axi_clk, arm_a9_hps:h2f_axi_clk, arm_a9_hps:h2f_lw_axi_clk, binaryscale:clk, greyparamter:clk, hps_vga_data1:clk, hps_vga_data2:clk, hwreset:clk, jtag_uart:clk, mm_interconnect_0:sdram_clk_sdram_clk_clk, mm_interconnect_1:sdram_clk_sdram_clk_clk, pio0:clk, pio_start:clk, rst_controller:clk, rst_controller_001:clk, sdram_to_hps_data1:clk, sdram_to_hps_data2:clk, sdramclock:clk, topedge:clk, vgabinary:clk, vgaclock:clk, vgaread:clk]
	wire          arm_a9_hps_h2f_axi_master_awvalid;                         // arm_a9_hps:h2f_AWVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awvalid
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;                          // arm_a9_hps:h2f_ARSIZE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arsize
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;                          // arm_a9_hps:h2f_ARLOCK -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arlock
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;                         // arm_a9_hps:h2f_AWCACHE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awcache
	wire          arm_a9_hps_h2f_axi_master_arready;                         // mm_interconnect_0:arm_a9_hps_h2f_axi_master_arready -> arm_a9_hps:h2f_ARREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;                            // arm_a9_hps:h2f_ARID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arid
	wire          arm_a9_hps_h2f_axi_master_rready;                          // arm_a9_hps:h2f_RREADY -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_rready
	wire          arm_a9_hps_h2f_axi_master_bready;                          // arm_a9_hps:h2f_BREADY -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_bready
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;                          // arm_a9_hps:h2f_AWSIZE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awsize
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;                          // arm_a9_hps:h2f_AWPROT -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awprot
	wire          arm_a9_hps_h2f_axi_master_arvalid;                         // arm_a9_hps:h2f_ARVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arvalid
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;                          // arm_a9_hps:h2f_ARPROT -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arprot
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;                             // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bid -> arm_a9_hps:h2f_BID
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;                           // arm_a9_hps:h2f_ARLEN -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arlen
	wire          arm_a9_hps_h2f_axi_master_awready;                         // mm_interconnect_0:arm_a9_hps_h2f_axi_master_awready -> arm_a9_hps:h2f_AWREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;                            // arm_a9_hps:h2f_AWID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awid
	wire          arm_a9_hps_h2f_axi_master_bvalid;                          // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bvalid -> arm_a9_hps:h2f_BVALID
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;                             // arm_a9_hps:h2f_WID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wid
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;                          // arm_a9_hps:h2f_AWLOCK -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;                         // arm_a9_hps:h2f_AWBURST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awburst
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;                           // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bresp -> arm_a9_hps:h2f_BRESP
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;                           // arm_a9_hps:h2f_WSTRB -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_rvalid;                          // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rvalid -> arm_a9_hps:h2f_RVALID
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;                           // arm_a9_hps:h2f_WDATA -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_wready;                          // mm_interconnect_0:arm_a9_hps_h2f_axi_master_wready -> arm_a9_hps:h2f_WREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;                         // arm_a9_hps:h2f_ARBURST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arburst
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;                           // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rdata -> arm_a9_hps:h2f_RDATA
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;                          // arm_a9_hps:h2f_ARADDR -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_araddr
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;                         // arm_a9_hps:h2f_ARCACHE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arcache
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;                           // arm_a9_hps:h2f_AWLEN -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awlen
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;                          // arm_a9_hps:h2f_AWADDR -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awaddr
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;                             // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rid -> arm_a9_hps:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_wvalid;                          // arm_a9_hps:h2f_WVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wvalid
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;                           // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rresp -> arm_a9_hps:h2f_RRESP
	wire          arm_a9_hps_h2f_axi_master_wlast;                           // arm_a9_hps:h2f_WLAST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wlast
	wire          arm_a9_hps_h2f_axi_master_rlast;                           // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rlast -> arm_a9_hps:h2f_RLAST
	wire   [31:0] mm_interconnect_0_onchip_sram_s1_writedata;                // mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire   [11:0] mm_interconnect_0_onchip_sram_s1_address;                  // mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire          mm_interconnect_0_onchip_sram_s1_chipselect;               // mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire          mm_interconnect_0_onchip_sram_s1_clken;                    // mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire          mm_interconnect_0_onchip_sram_s1_write;                    // mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire   [31:0] mm_interconnect_0_onchip_sram_s1_readdata;                 // Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	wire    [3:0] mm_interconnect_0_onchip_sram_s1_byteenable;               // mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire          arm_a9_hps_h2f_lw_axi_master_awvalid;                      // arm_a9_hps:h2f_lw_AWVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awvalid
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                       // arm_a9_hps:h2f_lw_ARSIZE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arsize
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                       // arm_a9_hps:h2f_lw_ARLOCK -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arlock
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                      // arm_a9_hps:h2f_lw_AWCACHE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awcache
	wire          arm_a9_hps_h2f_lw_axi_master_arready;                      // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arready -> arm_a9_hps:h2f_lw_ARREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                         // arm_a9_hps:h2f_lw_ARID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arid
	wire          arm_a9_hps_h2f_lw_axi_master_rready;                       // arm_a9_hps:h2f_lw_RREADY -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rready
	wire          arm_a9_hps_h2f_lw_axi_master_bready;                       // arm_a9_hps:h2f_lw_BREADY -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bready
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                       // arm_a9_hps:h2f_lw_AWSIZE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awsize
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                       // arm_a9_hps:h2f_lw_AWPROT -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awprot
	wire          arm_a9_hps_h2f_lw_axi_master_arvalid;                      // arm_a9_hps:h2f_lw_ARVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arvalid
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                       // arm_a9_hps:h2f_lw_ARPROT -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arprot
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                          // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bid -> arm_a9_hps:h2f_lw_BID
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                        // arm_a9_hps:h2f_lw_ARLEN -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arlen
	wire          arm_a9_hps_h2f_lw_axi_master_awready;                      // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awready -> arm_a9_hps:h2f_lw_AWREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                         // arm_a9_hps:h2f_lw_AWID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awid
	wire          arm_a9_hps_h2f_lw_axi_master_bvalid;                       // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bvalid -> arm_a9_hps:h2f_lw_BVALID
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                          // arm_a9_hps:h2f_lw_WID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                       // arm_a9_hps:h2f_lw_AWLOCK -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awlock
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                      // arm_a9_hps:h2f_lw_AWBURST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awburst
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                        // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bresp -> arm_a9_hps:h2f_lw_BRESP
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                        // arm_a9_hps:h2f_lw_WSTRB -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wstrb
	wire          arm_a9_hps_h2f_lw_axi_master_rvalid;                       // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rvalid -> arm_a9_hps:h2f_lw_RVALID
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                        // arm_a9_hps:h2f_lw_WDATA -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wdata
	wire          arm_a9_hps_h2f_lw_axi_master_wready;                       // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wready -> arm_a9_hps:h2f_lw_WREADY
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                      // arm_a9_hps:h2f_lw_ARBURST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arburst
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                        // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rdata -> arm_a9_hps:h2f_lw_RDATA
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                       // arm_a9_hps:h2f_lw_ARADDR -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_araddr
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                      // arm_a9_hps:h2f_lw_ARCACHE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arcache
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                        // arm_a9_hps:h2f_lw_AWLEN -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awlen
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                       // arm_a9_hps:h2f_lw_AWADDR -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awaddr
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                          // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rid -> arm_a9_hps:h2f_lw_RID
	wire          arm_a9_hps_h2f_lw_axi_master_wvalid;                       // arm_a9_hps:h2f_lw_WVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wvalid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                        // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rresp -> arm_a9_hps:h2f_lw_RRESP
	wire          arm_a9_hps_h2f_lw_axi_master_wlast;                        // arm_a9_hps:h2f_lw_WLAST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wlast
	wire          arm_a9_hps_h2f_lw_axi_master_rlast;                        // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rlast -> arm_a9_hps:h2f_lw_RLAST
	wire   [31:0] mm_interconnect_1_fifowe_s1_writedata;                     // mm_interconnect_1:FIFOWe_s1_writedata -> FIFOWe:writedata
	wire    [1:0] mm_interconnect_1_fifowe_s1_address;                       // mm_interconnect_1:FIFOWe_s1_address -> FIFOWe:address
	wire          mm_interconnect_1_fifowe_s1_chipselect;                    // mm_interconnect_1:FIFOWe_s1_chipselect -> FIFOWe:chipselect
	wire          mm_interconnect_1_fifowe_s1_write;                         // mm_interconnect_1:FIFOWe_s1_write -> FIFOWe:write_n
	wire   [31:0] mm_interconnect_1_fifowe_s1_readdata;                      // FIFOWe:readdata -> mm_interconnect_1:FIFOWe_s1_readdata
	wire   [31:0] mm_interconnect_1_hwreset_s1_writedata;                    // mm_interconnect_1:hwreset_s1_writedata -> hwreset:writedata
	wire    [1:0] mm_interconnect_1_hwreset_s1_address;                      // mm_interconnect_1:hwreset_s1_address -> hwreset:address
	wire          mm_interconnect_1_hwreset_s1_chipselect;                   // mm_interconnect_1:hwreset_s1_chipselect -> hwreset:chipselect
	wire          mm_interconnect_1_hwreset_s1_write;                        // mm_interconnect_1:hwreset_s1_write -> hwreset:write_n
	wire   [31:0] mm_interconnect_1_hwreset_s1_readdata;                     // hwreset:readdata -> mm_interconnect_1:hwreset_s1_readdata
	wire    [1:0] mm_interconnect_1_topedge_s1_address;                      // mm_interconnect_1:topedge_s1_address -> topedge:address
	wire   [31:0] mm_interconnect_1_topedge_s1_readdata;                     // topedge:readdata -> mm_interconnect_1:topedge_s1_readdata
	wire   [31:0] mm_interconnect_1_sdramclock_s1_writedata;                 // mm_interconnect_1:sdramclock_s1_writedata -> sdramclock:writedata
	wire    [1:0] mm_interconnect_1_sdramclock_s1_address;                   // mm_interconnect_1:sdramclock_s1_address -> sdramclock:address
	wire          mm_interconnect_1_sdramclock_s1_chipselect;                // mm_interconnect_1:sdramclock_s1_chipselect -> sdramclock:chipselect
	wire          mm_interconnect_1_sdramclock_s1_write;                     // mm_interconnect_1:sdramclock_s1_write -> sdramclock:write_n
	wire   [31:0] mm_interconnect_1_sdramclock_s1_readdata;                  // sdramclock:readdata -> mm_interconnect_1:sdramclock_s1_readdata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire    [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire   [31:0] mm_interconnect_1_greyparamter_s1_writedata;               // mm_interconnect_1:greyparamter_s1_writedata -> greyparamter:writedata
	wire    [1:0] mm_interconnect_1_greyparamter_s1_address;                 // mm_interconnect_1:greyparamter_s1_address -> greyparamter:address
	wire          mm_interconnect_1_greyparamter_s1_chipselect;              // mm_interconnect_1:greyparamter_s1_chipselect -> greyparamter:chipselect
	wire          mm_interconnect_1_greyparamter_s1_write;                   // mm_interconnect_1:greyparamter_s1_write -> greyparamter:write_n
	wire   [31:0] mm_interconnect_1_greyparamter_s1_readdata;                // greyparamter:readdata -> mm_interconnect_1:greyparamter_s1_readdata
	wire    [1:0] mm_interconnect_1_sdram_to_hps_data2_s1_address;           // mm_interconnect_1:sdram_to_hps_data2_s1_address -> sdram_to_hps_data2:address
	wire   [31:0] mm_interconnect_1_sdram_to_hps_data2_s1_readdata;          // sdram_to_hps_data2:readdata -> mm_interconnect_1:sdram_to_hps_data2_s1_readdata
	wire   [31:0] mm_interconnect_1_sdram_start_s1_writedata;                // mm_interconnect_1:Sdram_start_s1_writedata -> Sdram_start:writedata
	wire    [1:0] mm_interconnect_1_sdram_start_s1_address;                  // mm_interconnect_1:Sdram_start_s1_address -> Sdram_start:address
	wire          mm_interconnect_1_sdram_start_s1_chipselect;               // mm_interconnect_1:Sdram_start_s1_chipselect -> Sdram_start:chipselect
	wire          mm_interconnect_1_sdram_start_s1_write;                    // mm_interconnect_1:Sdram_start_s1_write -> Sdram_start:write_n
	wire   [31:0] mm_interconnect_1_sdram_start_s1_readdata;                 // Sdram_start:readdata -> mm_interconnect_1:Sdram_start_s1_readdata
	wire    [1:0] mm_interconnect_1_lval_s1_address;                         // mm_interconnect_1:Lval_s1_address -> Lval:address
	wire   [31:0] mm_interconnect_1_lval_s1_readdata;                        // Lval:readdata -> mm_interconnect_1:Lval_s1_readdata
	wire    [1:0] mm_interconnect_1_vgaclock_s1_address;                     // mm_interconnect_1:vgaclock_s1_address -> vgaclock:address
	wire   [31:0] mm_interconnect_1_vgaclock_s1_readdata;                    // vgaclock:readdata -> mm_interconnect_1:vgaclock_s1_readdata
	wire   [31:0] mm_interconnect_1_hps_vga_data1_s1_writedata;              // mm_interconnect_1:hps_vga_data1_s1_writedata -> hps_vga_data1:writedata
	wire    [1:0] mm_interconnect_1_hps_vga_data1_s1_address;                // mm_interconnect_1:hps_vga_data1_s1_address -> hps_vga_data1:address
	wire          mm_interconnect_1_hps_vga_data1_s1_chipselect;             // mm_interconnect_1:hps_vga_data1_s1_chipselect -> hps_vga_data1:chipselect
	wire          mm_interconnect_1_hps_vga_data1_s1_write;                  // mm_interconnect_1:hps_vga_data1_s1_write -> hps_vga_data1:write_n
	wire   [31:0] mm_interconnect_1_hps_vga_data1_s1_readdata;               // hps_vga_data1:readdata -> mm_interconnect_1:hps_vga_data1_s1_readdata
	wire   [31:0] mm_interconnect_1_hps_vga_data2_s1_writedata;              // mm_interconnect_1:hps_vga_data2_s1_writedata -> hps_vga_data2:writedata
	wire    [1:0] mm_interconnect_1_hps_vga_data2_s1_address;                // mm_interconnect_1:hps_vga_data2_s1_address -> hps_vga_data2:address
	wire          mm_interconnect_1_hps_vga_data2_s1_chipselect;             // mm_interconnect_1:hps_vga_data2_s1_chipselect -> hps_vga_data2:chipselect
	wire          mm_interconnect_1_hps_vga_data2_s1_write;                  // mm_interconnect_1:hps_vga_data2_s1_write -> hps_vga_data2:write_n
	wire   [31:0] mm_interconnect_1_hps_vga_data2_s1_readdata;               // hps_vga_data2:readdata -> mm_interconnect_1:hps_vga_data2_s1_readdata
	wire    [1:0] mm_interconnect_1_vgaread_s1_address;                      // mm_interconnect_1:vgaread_s1_address -> vgaread:address
	wire   [31:0] mm_interconnect_1_vgaread_s1_readdata;                     // vgaread:readdata -> mm_interconnect_1:vgaread_s1_readdata
	wire    [1:0] mm_interconnect_1_binaryscale_s1_address;                  // mm_interconnect_1:binaryscale_s1_address -> binaryscale:address
	wire   [31:0] mm_interconnect_1_binaryscale_s1_readdata;                 // binaryscale:readdata -> mm_interconnect_1:binaryscale_s1_readdata
	wire   [31:0] mm_interconnect_1_pio_start_s1_writedata;                  // mm_interconnect_1:pio_start_s1_writedata -> pio_start:writedata
	wire    [1:0] mm_interconnect_1_pio_start_s1_address;                    // mm_interconnect_1:pio_start_s1_address -> pio_start:address
	wire          mm_interconnect_1_pio_start_s1_chipselect;                 // mm_interconnect_1:pio_start_s1_chipselect -> pio_start:chipselect
	wire          mm_interconnect_1_pio_start_s1_write;                      // mm_interconnect_1:pio_start_s1_write -> pio_start:write_n
	wire   [31:0] mm_interconnect_1_pio_start_s1_readdata;                   // pio_start:readdata -> mm_interconnect_1:pio_start_s1_readdata
	wire   [31:0] mm_interconnect_1_vgabinary_s1_writedata;                  // mm_interconnect_1:vgabinary_s1_writedata -> vgabinary:writedata
	wire    [1:0] mm_interconnect_1_vgabinary_s1_address;                    // mm_interconnect_1:vgabinary_s1_address -> vgabinary:address
	wire          mm_interconnect_1_vgabinary_s1_chipselect;                 // mm_interconnect_1:vgabinary_s1_chipselect -> vgabinary:chipselect
	wire          mm_interconnect_1_vgabinary_s1_write;                      // mm_interconnect_1:vgabinary_s1_write -> vgabinary:write_n
	wire   [31:0] mm_interconnect_1_vgabinary_s1_readdata;                   // vgabinary:readdata -> mm_interconnect_1:vgabinary_s1_readdata
	wire   [31:0] mm_interconnect_1_pio0_s1_writedata;                       // mm_interconnect_1:pio0_s1_writedata -> pio0:writedata
	wire    [1:0] mm_interconnect_1_pio0_s1_address;                         // mm_interconnect_1:pio0_s1_address -> pio0:address
	wire          mm_interconnect_1_pio0_s1_chipselect;                      // mm_interconnect_1:pio0_s1_chipselect -> pio0:chipselect
	wire          mm_interconnect_1_pio0_s1_write;                           // mm_interconnect_1:pio0_s1_write -> pio0:write_n
	wire   [31:0] mm_interconnect_1_pio0_s1_readdata;                        // pio0:readdata -> mm_interconnect_1:pio0_s1_readdata
	wire    [1:0] mm_interconnect_1_sdram_to_hps_data1_s1_address;           // mm_interconnect_1:sdram_to_hps_data1_s1_address -> sdram_to_hps_data1:address
	wire   [31:0] mm_interconnect_1_sdram_to_hps_data1_s1_readdata;          // sdram_to_hps_data1:readdata -> mm_interconnect_1:sdram_to_hps_data1_s1_readdata
	wire          irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                                   // irq_mapper:sender_irq -> arm_a9_hps:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                                   // irq_mapper_001:sender_irq -> arm_a9_hps:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [FIFOWe:reset_n, Lval:reset_n, Onchip_SRAM:reset, Sdram_start:reset_n, binaryscale:reset_n, greyparamter:reset_n, hps_vga_data1:reset_n, hps_vga_data2:reset_n, hwreset:reset_n, jtag_uart:rst_n, mm_interconnect_0:Onchip_SRAM_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:pio0_reset_reset_bridge_in_reset_reset, pio0:reset_n, pio_start:reset_n, rst_translator:in_reset, sdram_to_hps_data1:reset_n, sdram_to_hps_data2:reset_n, sdramclock:reset_n, topedge:reset_n, vgabinary:reset_n, vgaclock:reset_n, vgaread:reset_n]
	wire          rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire          arm_a9_hps_h2f_reset_reset;                                // arm_a9_hps:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire          sdram_clk_reset_source_reset;                              // sdram_clk:reset_source_reset -> rst_controller:reset_in1
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_0:arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	mysystem_arm_a9_hps #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a          (memory_mem_a),                         //            memory.mem_a
		.mem_ba         (memory_mem_ba),                        //                  .mem_ba
		.mem_ck         (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n       (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke        (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n       (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n       (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq         (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs        (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt        (memory_mem_odt),                       //                  .mem_odt
		.mem_dm         (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin      (memory_oct_rzqin),                     //                  .oct_rzqin
		.h2f_rst_n      (arm_a9_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk    (sdram_clk_sdram_clk_clk),              //     h2f_axi_clock.clk
		.h2f_AWID       (arm_a9_hps_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR     (arm_a9_hps_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN      (arm_a9_hps_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE     (arm_a9_hps_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST    (arm_a9_hps_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK     (arm_a9_hps_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE    (arm_a9_hps_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT     (arm_a9_hps_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID    (arm_a9_hps_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY    (arm_a9_hps_h2f_axi_master_awready),    //                  .awready
		.h2f_WID        (arm_a9_hps_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA      (arm_a9_hps_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB      (arm_a9_hps_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST      (arm_a9_hps_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID     (arm_a9_hps_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY     (arm_a9_hps_h2f_axi_master_wready),     //                  .wready
		.h2f_BID        (arm_a9_hps_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP      (arm_a9_hps_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID     (arm_a9_hps_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY     (arm_a9_hps_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID       (arm_a9_hps_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR     (arm_a9_hps_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN      (arm_a9_hps_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE     (arm_a9_hps_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST    (arm_a9_hps_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK     (arm_a9_hps_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE    (arm_a9_hps_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT     (arm_a9_hps_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID    (arm_a9_hps_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY    (arm_a9_hps_h2f_axi_master_arready),    //                  .arready
		.h2f_RID        (arm_a9_hps_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA      (arm_a9_hps_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP      (arm_a9_hps_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST      (arm_a9_hps_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID     (arm_a9_hps_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY     (arm_a9_hps_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk    (sdram_clk_sdram_clk_clk),              //     f2h_axi_clock.clk
		.f2h_AWID       (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR     (),                                     //                  .awaddr
		.f2h_AWLEN      (),                                     //                  .awlen
		.f2h_AWSIZE     (),                                     //                  .awsize
		.f2h_AWBURST    (),                                     //                  .awburst
		.f2h_AWLOCK     (),                                     //                  .awlock
		.f2h_AWCACHE    (),                                     //                  .awcache
		.f2h_AWPROT     (),                                     //                  .awprot
		.f2h_AWVALID    (),                                     //                  .awvalid
		.f2h_AWREADY    (),                                     //                  .awready
		.f2h_AWUSER     (),                                     //                  .awuser
		.f2h_WID        (),                                     //                  .wid
		.f2h_WDATA      (),                                     //                  .wdata
		.f2h_WSTRB      (),                                     //                  .wstrb
		.f2h_WLAST      (),                                     //                  .wlast
		.f2h_WVALID     (),                                     //                  .wvalid
		.f2h_WREADY     (),                                     //                  .wready
		.f2h_BID        (),                                     //                  .bid
		.f2h_BRESP      (),                                     //                  .bresp
		.f2h_BVALID     (),                                     //                  .bvalid
		.f2h_BREADY     (),                                     //                  .bready
		.f2h_ARID       (),                                     //                  .arid
		.f2h_ARADDR     (),                                     //                  .araddr
		.f2h_ARLEN      (),                                     //                  .arlen
		.f2h_ARSIZE     (),                                     //                  .arsize
		.f2h_ARBURST    (),                                     //                  .arburst
		.f2h_ARLOCK     (),                                     //                  .arlock
		.f2h_ARCACHE    (),                                     //                  .arcache
		.f2h_ARPROT     (),                                     //                  .arprot
		.f2h_ARVALID    (),                                     //                  .arvalid
		.f2h_ARREADY    (),                                     //                  .arready
		.f2h_ARUSER     (),                                     //                  .aruser
		.f2h_RID        (),                                     //                  .rid
		.f2h_RDATA      (),                                     //                  .rdata
		.f2h_RRESP      (),                                     //                  .rresp
		.f2h_RLAST      (),                                     //                  .rlast
		.f2h_RVALID     (),                                     //                  .rvalid
		.f2h_RREADY     (),                                     //                  .rready
		.h2f_lw_axi_clk (sdram_clk_sdram_clk_clk),              //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (arm_a9_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (arm_a9_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN   (arm_a9_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE  (arm_a9_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST (arm_a9_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK  (arm_a9_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE (arm_a9_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT  (arm_a9_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID (arm_a9_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY (arm_a9_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID     (arm_a9_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA   (arm_a9_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB   (arm_a9_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST   (arm_a9_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID  (arm_a9_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY  (arm_a9_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID     (arm_a9_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP   (arm_a9_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID  (arm_a9_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY  (arm_a9_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID    (arm_a9_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR  (arm_a9_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN   (arm_a9_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE  (arm_a9_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST (arm_a9_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK  (arm_a9_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE (arm_a9_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT  (arm_a9_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID (arm_a9_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY (arm_a9_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID     (arm_a9_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA   (arm_a9_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP   (arm_a9_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST   (arm_a9_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID  (arm_a9_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY  (arm_a9_hps_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0     (arm_a9_hps_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1     (arm_a9_hps_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	mysystem_pio0 pio0 (
		.clk        (sdram_clk_sdram_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_pio0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio0_s1_readdata),   //                    .readdata
		.out_port   (hps_read_export)                       // external_connection.export
	);

	mysystem_jtag_uart jtag_uart (
		.clk            (sdram_clk_sdram_clk_clk),                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	mysystem_Onchip_SRAM onchip_sram (
		.clk        (sdram_clk_sdram_clk_clk),                     //   clk1.clk
		.address    (mm_interconnect_0_onchip_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)           //       .reset_req
	);

	mysystem_system_pll_0 system_pll_0 (
		.refclk   (system_pll_0_refclk_clk),  //  refclk.clk
		.rst      (system_pll_0_reset_reset), //   reset.reset
		.outclk_0 (sdram_clk_clk),            // outclk0.clk
		.outclk_1 (dram_clk_clk),             // outclk1.clk
		.outclk_2 (d5m_clk_clk),              // outclk2.clk
		.outclk_3 (vga_clk_clk),              // outclk3.clk
		.locked   ()                          // (terminated)
	);

	mysystem_sdram_clk sdram_clk (
		.ref_clk_clk        (sdram_clk_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (sdram_clk_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (),                             //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_sdram_clk_clk),      //    sdram_clk.clk
		.reset_source_reset (sdram_clk_reset_source_reset)  // reset_source.reset
	);

	mysystem_sdram_to_hps_data2 sdram_to_hps_data2 (
		.clk      (sdram_clk_sdram_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_1_sdram_to_hps_data2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sdram_to_hps_data2_s1_readdata), //                    .readdata
		.in_port  (sdram_hps_data2_export)                            // external_connection.export
	);

	mysystem_sdram_to_hps_data2 sdram_to_hps_data1 (
		.clk      (sdram_clk_sdram_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_1_sdram_to_hps_data1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sdram_to_hps_data1_s1_readdata), //                    .readdata
		.in_port  (sdram_hps_data1_export)                            // external_connection.export
	);

	mysystem_pio0 pio_start (
		.clk        (sdram_clk_sdram_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_pio_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_start_s1_readdata),   //                    .readdata
		.out_port   (capture_start_export)                       // external_connection.export
	);

	mysystem_hps_vga_data1 hps_vga_data1 (
		.clk        (sdram_clk_sdram_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_1_hps_vga_data1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_hps_vga_data1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_hps_vga_data1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_hps_vga_data1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_hps_vga_data1_s1_readdata),   //                    .readdata
		.out_port   (hps_vga_data1_export)                           // external_connection.export
	);

	mysystem_hps_vga_data1 hps_vga_data2 (
		.clk        (sdram_clk_sdram_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_1_hps_vga_data2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_hps_vga_data2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_hps_vga_data2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_hps_vga_data2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_hps_vga_data2_s1_readdata),   //                    .readdata
		.out_port   (hps_vga_data2_export)                           // external_connection.export
	);

	mysystem_pio0 sdramclock (
		.clk        (sdram_clk_sdram_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_sdramclock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sdramclock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sdramclock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sdramclock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sdramclock_s1_readdata),   //                    .readdata
		.out_port   (sdramclock_export)                           // external_connection.export
	);

	mysystem_pio0 sdram_start (
		.clk        (sdram_clk_sdram_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_sdram_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sdram_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sdram_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sdram_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sdram_start_s1_readdata),   //                    .readdata
		.out_port   (sdram_start_export)                           // external_connection.export
	);

	mysystem_pio0 fifowe (
		.clk        (sdram_clk_sdram_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_fifowe_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_fifowe_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_fifowe_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_fifowe_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_fifowe_s1_readdata),   //                    .readdata
		.out_port   (fifowe_export)                           // external_connection.export
	);

	mysystem_binaryscale binaryscale (
		.clk      (sdram_clk_sdram_clk_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_binaryscale_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_binaryscale_s1_readdata), //                    .readdata
		.in_port  (binary_export)                              // external_connection.export
	);

	mysystem_greyparamter greyparamter (
		.clk        (sdram_clk_sdram_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_greyparamter_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_greyparamter_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_greyparamter_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_greyparamter_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_greyparamter_s1_readdata),   //                    .readdata
		.out_port   (greyparameter_export)                          // external_connection.export
	);

	mysystem_vgaclock vgaclock (
		.clk      (sdram_clk_sdram_clk_clk),                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_1_vgaclock_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_vgaclock_s1_readdata), //                    .readdata
		.in_port  (vgaclock_export)                         // external_connection.export
	);

	mysystem_pio0 vgabinary (
		.clk        (sdram_clk_sdram_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_vgabinary_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_vgabinary_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_vgabinary_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_vgabinary_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_vgabinary_s1_readdata),   //                    .readdata
		.out_port   (vgabinary_export)                           // external_connection.export
	);

	mysystem_vgaclock vgaread (
		.clk      (sdram_clk_sdram_clk_clk),               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_1_vgaread_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_vgaread_s1_readdata), //                    .readdata
		.in_port  (vgaread_export)                         // external_connection.export
	);

	mysystem_binaryscale topedge (
		.clk      (sdram_clk_sdram_clk_clk),               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_1_topedge_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_topedge_s1_readdata), //                    .readdata
		.in_port  (topedge_export)                         // external_connection.export
	);

	mysystem_pio0 hwreset (
		.clk        (sdram_clk_sdram_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_hwreset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_hwreset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_hwreset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_hwreset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_hwreset_s1_readdata),   //                    .readdata
		.out_port   (hwreset_export)                           // external_connection.export
	);

	mysystem_vgaclock lval (
		.clk      (sdram_clk_sdram_clk_clk),            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_1_lval_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_lval_s1_readdata), //                    .readdata
		.in_port  (lval_export)                         // external_connection.export
	);

	mysystem_mm_interconnect_0 mm_interconnect_0 (
		.arm_a9_hps_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),              //                                       arm_a9_hps_h2f_axi_master.awid
		.arm_a9_hps_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),            //                                                                .awaddr
		.arm_a9_hps_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),             //                                                                .awlen
		.arm_a9_hps_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),            //                                                                .awsize
		.arm_a9_hps_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),           //                                                                .awburst
		.arm_a9_hps_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),            //                                                                .awlock
		.arm_a9_hps_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),           //                                                                .awcache
		.arm_a9_hps_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),            //                                                                .awprot
		.arm_a9_hps_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),           //                                                                .awvalid
		.arm_a9_hps_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),           //                                                                .awready
		.arm_a9_hps_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),               //                                                                .wid
		.arm_a9_hps_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),             //                                                                .wdata
		.arm_a9_hps_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),             //                                                                .wstrb
		.arm_a9_hps_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),             //                                                                .wlast
		.arm_a9_hps_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),            //                                                                .wvalid
		.arm_a9_hps_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),            //                                                                .wready
		.arm_a9_hps_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),               //                                                                .bid
		.arm_a9_hps_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),             //                                                                .bresp
		.arm_a9_hps_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),            //                                                                .bvalid
		.arm_a9_hps_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),            //                                                                .bready
		.arm_a9_hps_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),              //                                                                .arid
		.arm_a9_hps_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),            //                                                                .araddr
		.arm_a9_hps_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),             //                                                                .arlen
		.arm_a9_hps_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),            //                                                                .arsize
		.arm_a9_hps_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),           //                                                                .arburst
		.arm_a9_hps_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),            //                                                                .arlock
		.arm_a9_hps_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),           //                                                                .arcache
		.arm_a9_hps_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),            //                                                                .arprot
		.arm_a9_hps_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),           //                                                                .arvalid
		.arm_a9_hps_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),           //                                                                .arready
		.arm_a9_hps_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),               //                                                                .rid
		.arm_a9_hps_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),             //                                                                .rdata
		.arm_a9_hps_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),             //                                                                .rresp
		.arm_a9_hps_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),             //                                                                .rlast
		.arm_a9_hps_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),            //                                                                .rvalid
		.arm_a9_hps_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),            //                                                                .rready
		.sdram_clk_sdram_clk_clk                                               (sdram_clk_sdram_clk_clk),                     //                                             sdram_clk_sdram_clk.clk
		.arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),          // arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Onchip_SRAM_reset1_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),              //                        Onchip_SRAM_reset1_reset_bridge_in_reset.reset
		.Onchip_SRAM_s1_address                                                (mm_interconnect_0_onchip_sram_s1_address),    //                                                  Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                                                  (mm_interconnect_0_onchip_sram_s1_write),      //                                                                .write
		.Onchip_SRAM_s1_readdata                                               (mm_interconnect_0_onchip_sram_s1_readdata),   //                                                                .readdata
		.Onchip_SRAM_s1_writedata                                              (mm_interconnect_0_onchip_sram_s1_writedata),  //                                                                .writedata
		.Onchip_SRAM_s1_byteenable                                             (mm_interconnect_0_onchip_sram_s1_byteenable), //                                                                .byteenable
		.Onchip_SRAM_s1_chipselect                                             (mm_interconnect_0_onchip_sram_s1_chipselect), //                                                                .chipselect
		.Onchip_SRAM_s1_clken                                                  (mm_interconnect_0_onchip_sram_s1_clken)       //                                                                .clken
	);

	mysystem_mm_interconnect_1 mm_interconnect_1 (
		.arm_a9_hps_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                         //                                       arm_a9_hps_h2f_lw_axi_master.awid
		.arm_a9_hps_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                       //                                                                   .awaddr
		.arm_a9_hps_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                        //                                                                   .awlen
		.arm_a9_hps_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                       //                                                                   .awsize
		.arm_a9_hps_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                      //                                                                   .awburst
		.arm_a9_hps_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                       //                                                                   .awlock
		.arm_a9_hps_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                      //                                                                   .awcache
		.arm_a9_hps_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                       //                                                                   .awprot
		.arm_a9_hps_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                      //                                                                   .awvalid
		.arm_a9_hps_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                      //                                                                   .awready
		.arm_a9_hps_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                          //                                                                   .wid
		.arm_a9_hps_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                        //                                                                   .wdata
		.arm_a9_hps_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                        //                                                                   .wstrb
		.arm_a9_hps_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                        //                                                                   .wlast
		.arm_a9_hps_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                       //                                                                   .wvalid
		.arm_a9_hps_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                       //                                                                   .wready
		.arm_a9_hps_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                          //                                                                   .bid
		.arm_a9_hps_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                        //                                                                   .bresp
		.arm_a9_hps_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                       //                                                                   .bvalid
		.arm_a9_hps_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                       //                                                                   .bready
		.arm_a9_hps_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                         //                                                                   .arid
		.arm_a9_hps_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                       //                                                                   .araddr
		.arm_a9_hps_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                        //                                                                   .arlen
		.arm_a9_hps_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                       //                                                                   .arsize
		.arm_a9_hps_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                      //                                                                   .arburst
		.arm_a9_hps_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                       //                                                                   .arlock
		.arm_a9_hps_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                      //                                                                   .arcache
		.arm_a9_hps_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                       //                                                                   .arprot
		.arm_a9_hps_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                      //                                                                   .arvalid
		.arm_a9_hps_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                      //                                                                   .arready
		.arm_a9_hps_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                          //                                                                   .rid
		.arm_a9_hps_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                        //                                                                   .rdata
		.arm_a9_hps_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                        //                                                                   .rresp
		.arm_a9_hps_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                        //                                                                   .rlast
		.arm_a9_hps_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                       //                                                                   .rvalid
		.arm_a9_hps_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                       //                                                                   .rready
		.sdram_clk_sdram_clk_clk                                                  (sdram_clk_sdram_clk_clk),                                   //                                                sdram_clk_sdram_clk.clk
		.arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio0_reset_reset_bridge_in_reset_reset                                   (rst_controller_reset_out_reset),                            //                                   pio0_reset_reset_bridge_in_reset.reset
		.binaryscale_s1_address                                                   (mm_interconnect_1_binaryscale_s1_address),                  //                                                     binaryscale_s1.address
		.binaryscale_s1_readdata                                                  (mm_interconnect_1_binaryscale_s1_readdata),                 //                                                                   .readdata
		.FIFOWe_s1_address                                                        (mm_interconnect_1_fifowe_s1_address),                       //                                                          FIFOWe_s1.address
		.FIFOWe_s1_write                                                          (mm_interconnect_1_fifowe_s1_write),                         //                                                                   .write
		.FIFOWe_s1_readdata                                                       (mm_interconnect_1_fifowe_s1_readdata),                      //                                                                   .readdata
		.FIFOWe_s1_writedata                                                      (mm_interconnect_1_fifowe_s1_writedata),                     //                                                                   .writedata
		.FIFOWe_s1_chipselect                                                     (mm_interconnect_1_fifowe_s1_chipselect),                    //                                                                   .chipselect
		.greyparamter_s1_address                                                  (mm_interconnect_1_greyparamter_s1_address),                 //                                                    greyparamter_s1.address
		.greyparamter_s1_write                                                    (mm_interconnect_1_greyparamter_s1_write),                   //                                                                   .write
		.greyparamter_s1_readdata                                                 (mm_interconnect_1_greyparamter_s1_readdata),                //                                                                   .readdata
		.greyparamter_s1_writedata                                                (mm_interconnect_1_greyparamter_s1_writedata),               //                                                                   .writedata
		.greyparamter_s1_chipselect                                               (mm_interconnect_1_greyparamter_s1_chipselect),              //                                                                   .chipselect
		.hps_vga_data1_s1_address                                                 (mm_interconnect_1_hps_vga_data1_s1_address),                //                                                   hps_vga_data1_s1.address
		.hps_vga_data1_s1_write                                                   (mm_interconnect_1_hps_vga_data1_s1_write),                  //                                                                   .write
		.hps_vga_data1_s1_readdata                                                (mm_interconnect_1_hps_vga_data1_s1_readdata),               //                                                                   .readdata
		.hps_vga_data1_s1_writedata                                               (mm_interconnect_1_hps_vga_data1_s1_writedata),              //                                                                   .writedata
		.hps_vga_data1_s1_chipselect                                              (mm_interconnect_1_hps_vga_data1_s1_chipselect),             //                                                                   .chipselect
		.hps_vga_data2_s1_address                                                 (mm_interconnect_1_hps_vga_data2_s1_address),                //                                                   hps_vga_data2_s1.address
		.hps_vga_data2_s1_write                                                   (mm_interconnect_1_hps_vga_data2_s1_write),                  //                                                                   .write
		.hps_vga_data2_s1_readdata                                                (mm_interconnect_1_hps_vga_data2_s1_readdata),               //                                                                   .readdata
		.hps_vga_data2_s1_writedata                                               (mm_interconnect_1_hps_vga_data2_s1_writedata),              //                                                                   .writedata
		.hps_vga_data2_s1_chipselect                                              (mm_interconnect_1_hps_vga_data2_s1_chipselect),             //                                                                   .chipselect
		.hwreset_s1_address                                                       (mm_interconnect_1_hwreset_s1_address),                      //                                                         hwreset_s1.address
		.hwreset_s1_write                                                         (mm_interconnect_1_hwreset_s1_write),                        //                                                                   .write
		.hwreset_s1_readdata                                                      (mm_interconnect_1_hwreset_s1_readdata),                     //                                                                   .readdata
		.hwreset_s1_writedata                                                     (mm_interconnect_1_hwreset_s1_writedata),                    //                                                                   .writedata
		.hwreset_s1_chipselect                                                    (mm_interconnect_1_hwreset_s1_chipselect),                   //                                                                   .chipselect
		.jtag_uart_avalon_jtag_slave_address                                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                                   .write
		.jtag_uart_avalon_jtag_slave_read                                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                                   .chipselect
		.Lval_s1_address                                                          (mm_interconnect_1_lval_s1_address),                         //                                                            Lval_s1.address
		.Lval_s1_readdata                                                         (mm_interconnect_1_lval_s1_readdata),                        //                                                                   .readdata
		.pio0_s1_address                                                          (mm_interconnect_1_pio0_s1_address),                         //                                                            pio0_s1.address
		.pio0_s1_write                                                            (mm_interconnect_1_pio0_s1_write),                           //                                                                   .write
		.pio0_s1_readdata                                                         (mm_interconnect_1_pio0_s1_readdata),                        //                                                                   .readdata
		.pio0_s1_writedata                                                        (mm_interconnect_1_pio0_s1_writedata),                       //                                                                   .writedata
		.pio0_s1_chipselect                                                       (mm_interconnect_1_pio0_s1_chipselect),                      //                                                                   .chipselect
		.pio_start_s1_address                                                     (mm_interconnect_1_pio_start_s1_address),                    //                                                       pio_start_s1.address
		.pio_start_s1_write                                                       (mm_interconnect_1_pio_start_s1_write),                      //                                                                   .write
		.pio_start_s1_readdata                                                    (mm_interconnect_1_pio_start_s1_readdata),                   //                                                                   .readdata
		.pio_start_s1_writedata                                                   (mm_interconnect_1_pio_start_s1_writedata),                  //                                                                   .writedata
		.pio_start_s1_chipselect                                                  (mm_interconnect_1_pio_start_s1_chipselect),                 //                                                                   .chipselect
		.Sdram_start_s1_address                                                   (mm_interconnect_1_sdram_start_s1_address),                  //                                                     Sdram_start_s1.address
		.Sdram_start_s1_write                                                     (mm_interconnect_1_sdram_start_s1_write),                    //                                                                   .write
		.Sdram_start_s1_readdata                                                  (mm_interconnect_1_sdram_start_s1_readdata),                 //                                                                   .readdata
		.Sdram_start_s1_writedata                                                 (mm_interconnect_1_sdram_start_s1_writedata),                //                                                                   .writedata
		.Sdram_start_s1_chipselect                                                (mm_interconnect_1_sdram_start_s1_chipselect),               //                                                                   .chipselect
		.sdram_to_hps_data1_s1_address                                            (mm_interconnect_1_sdram_to_hps_data1_s1_address),           //                                              sdram_to_hps_data1_s1.address
		.sdram_to_hps_data1_s1_readdata                                           (mm_interconnect_1_sdram_to_hps_data1_s1_readdata),          //                                                                   .readdata
		.sdram_to_hps_data2_s1_address                                            (mm_interconnect_1_sdram_to_hps_data2_s1_address),           //                                              sdram_to_hps_data2_s1.address
		.sdram_to_hps_data2_s1_readdata                                           (mm_interconnect_1_sdram_to_hps_data2_s1_readdata),          //                                                                   .readdata
		.sdramclock_s1_address                                                    (mm_interconnect_1_sdramclock_s1_address),                   //                                                      sdramclock_s1.address
		.sdramclock_s1_write                                                      (mm_interconnect_1_sdramclock_s1_write),                     //                                                                   .write
		.sdramclock_s1_readdata                                                   (mm_interconnect_1_sdramclock_s1_readdata),                  //                                                                   .readdata
		.sdramclock_s1_writedata                                                  (mm_interconnect_1_sdramclock_s1_writedata),                 //                                                                   .writedata
		.sdramclock_s1_chipselect                                                 (mm_interconnect_1_sdramclock_s1_chipselect),                //                                                                   .chipselect
		.topedge_s1_address                                                       (mm_interconnect_1_topedge_s1_address),                      //                                                         topedge_s1.address
		.topedge_s1_readdata                                                      (mm_interconnect_1_topedge_s1_readdata),                     //                                                                   .readdata
		.vgabinary_s1_address                                                     (mm_interconnect_1_vgabinary_s1_address),                    //                                                       vgabinary_s1.address
		.vgabinary_s1_write                                                       (mm_interconnect_1_vgabinary_s1_write),                      //                                                                   .write
		.vgabinary_s1_readdata                                                    (mm_interconnect_1_vgabinary_s1_readdata),                   //                                                                   .readdata
		.vgabinary_s1_writedata                                                   (mm_interconnect_1_vgabinary_s1_writedata),                  //                                                                   .writedata
		.vgabinary_s1_chipselect                                                  (mm_interconnect_1_vgabinary_s1_chipselect),                 //                                                                   .chipselect
		.vgaclock_s1_address                                                      (mm_interconnect_1_vgaclock_s1_address),                     //                                                        vgaclock_s1.address
		.vgaclock_s1_readdata                                                     (mm_interconnect_1_vgaclock_s1_readdata),                    //                                                                   .readdata
		.vgaread_s1_address                                                       (mm_interconnect_1_vgaread_s1_address),                      //                                                         vgaread_s1.address
		.vgaread_s1_readdata                                                      (mm_interconnect_1_vgaread_s1_readdata)                      //                                                                   .readdata
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	mysystem_irq_mapper_001 irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (sdram_clk_reset_source_reset),       // reset_in1.reset
		.clk            (sdram_clk_sdram_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (sdram_clk_sdram_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
